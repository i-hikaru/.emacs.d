-------------------------------------------------------------------------------
-- file name:      
-- author:         hikaru
--
-- create date:    
-- module name:    
-- project name:   
-- target devices: 
-- tool versions:  
-- description:    
-- dependencies:   
--
-- revision:       
-- comments:       
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--library unisim;
--use unisim.vcomponents.all;
