--------------------------------------------------------------------------------
-- file name: 
-- author:
--
-- create date: 
-- module name: 
-- project name: 
-- target devices: 
-- versions: 
-- description: 
-- dependencies: 
--
-- revision: 
-- comments: 
--
--------------------------------------------------------------------------------
